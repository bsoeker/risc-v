library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity rom is
    generic (
        addr_width  : integer := 12;  -- 2^10 = 1KB
        data_width  : integer := 32 
    );
    port (
        instr_addr : in  std_logic_vector(addr_width - 1 downto 0); -- Byte address (PC)
        instr_data : out std_logic_vector(data_width - 1 downto 0);  -- Full 32-bit instruction
        data_addr : in  std_logic_vector(addr_width - 1 downto 0); -- Byte address (ALU)
        data_data : out std_logic_vector(data_width - 1 downto 0)  -- Full 32-bit data

    );
end rom;

architecture rom_arch of rom is

    -- Byte-addressable ROM: Each address holds 1 byte
    type rom_type is array (0 to 2**addr_width - 1) of std_logic_vector(7 downto 0);
    signal rom_array : rom_type := (
    0 => x"17",
    1 => x"11",
    2 => x"00",
    3 => x"10",
    4 => x"13",
    5 => x"01",
    6 => x"01",
    7 => x"00",
    8 => x"13",
    9 => x"05",
    10 => x"40",
    11 => x"0E",
    12 => x"97",
    13 => x"05",
    14 => x"00",
    15 => x"10",
    16 => x"93",
    17 => x"85",
    18 => x"45",
    19 => x"FF",
    20 => x"17",
    21 => x"06",
    22 => x"00",
    23 => x"10",
    24 => x"13",
    25 => x"06",
    26 => x"26",
    27 => x"FF",
    28 => x"63",
    29 => x"8C",
    30 => x"C5",
    31 => x"00",
    32 => x"83",
    33 => x"42",
    34 => x"05",
    35 => x"00",
    36 => x"23",
    37 => x"80",
    38 => x"55",
    39 => x"00",
    40 => x"13",
    41 => x"05",
    42 => x"15",
    43 => x"00",
    44 => x"93",
    45 => x"85",
    46 => x"15",
    47 => x"00",
    48 => x"6F",
    49 => x"F0",
    50 => x"DF",
    51 => x"FE",
    52 => x"17",
    53 => x"05",
    54 => x"00",
    55 => x"10",
    56 => x"13",
    57 => x"05",
    58 => x"25",
    59 => x"FD",
    60 => x"97",
    61 => x"05",
    62 => x"00",
    63 => x"10",
    64 => x"93",
    65 => x"85",
    66 => x"A5",
    67 => x"FC",
    68 => x"63",
    69 => x"08",
    70 => x"B5",
    71 => x"00",
    72 => x"23",
    73 => x"20",
    74 => x"05",
    75 => x"00",
    76 => x"13",
    77 => x"05",
    78 => x"45",
    79 => x"00",
    80 => x"6F",
    81 => x"F0",
    82 => x"5F",
    83 => x"FF",
    84 => x"EF",
    85 => x"00",
    86 => x"40",
    87 => x"05",
    88 => x"6F",
    89 => x"00",
    90 => x"00",
    91 => x"00",
    92 => x"13",
    93 => x"01",
    94 => x"01",
    95 => x"FE",
    96 => x"23",
    97 => x"2E",
    98 => x"11",
    99 => x"00",
    100 => x"23",
    101 => x"2C",
    102 => x"81",
    103 => x"00",
    104 => x"13",
    105 => x"04",
    106 => x"01",
    107 => x"02",
    108 => x"23",
    109 => x"26",
    110 => x"04",
    111 => x"FE",
    112 => x"6F",
    113 => x"00",
    114 => x"00",
    115 => x"01",
    116 => x"83",
    117 => x"27",
    118 => x"C4",
    119 => x"FE",
    120 => x"93",
    121 => x"87",
    122 => x"17",
    123 => x"00",
    124 => x"23",
    125 => x"26",
    126 => x"F4",
    127 => x"FE",
    128 => x"03",
    129 => x"27",
    130 => x"C4",
    131 => x"FE",
    132 => x"B7",
    133 => x"47",
    134 => x"0F",
    135 => x"00",
    136 => x"93",
    137 => x"87",
    138 => x"F7",
    139 => x"23",
    140 => x"E3",
    141 => x"D4",
    142 => x"E7",
    143 => x"FE",
    144 => x"13",
    145 => x"00",
    146 => x"00",
    147 => x"00",
    148 => x"13",
    149 => x"00",
    150 => x"00",
    151 => x"00",
    152 => x"83",
    153 => x"20",
    154 => x"C1",
    155 => x"01",
    156 => x"03",
    157 => x"24",
    158 => x"81",
    159 => x"01",
    160 => x"13",
    161 => x"01",
    162 => x"01",
    163 => x"02",
    164 => x"67",
    165 => x"80",
    166 => x"00",
    167 => x"00",
    168 => x"13",
    169 => x"01",
    170 => x"01",
    171 => x"FF",
    172 => x"23",
    173 => x"26",
    174 => x"11",
    175 => x"00",
    176 => x"23",
    177 => x"24",
    178 => x"81",
    179 => x"00",
    180 => x"13",
    181 => x"04",
    182 => x"01",
    183 => x"01",
    184 => x"B7",
    185 => x"07",
    186 => x"00",
    187 => x"10",
    188 => x"93",
    189 => x"87",
    190 => x"07",
    191 => x"00",
    192 => x"03",
    193 => x"C7",
    194 => x"07",
    195 => x"00",
    196 => x"B7",
    197 => x"07",
    198 => x"00",
    199 => x"20",
    200 => x"23",
    201 => x"A0",
    202 => x"E7",
    203 => x"00",
    204 => x"93",
    205 => x"07",
    206 => x"00",
    207 => x"00",
    208 => x"13",
    209 => x"85",
    210 => x"07",
    211 => x"00",
    212 => x"83",
    213 => x"20",
    214 => x"C1",
    215 => x"00",
    216 => x"03",
    217 => x"24",
    218 => x"81",
    219 => x"00",
    220 => x"13",
    221 => x"01",
    222 => x"01",
    223 => x"01",
    224 => x"67",
    225 => x"80",
    226 => x"00",
    227 => x"00",
    228 => x"48",
    229 => x"65",
    230 => x"6C",
    231 => x"6C",
    232 => x"6F",
    233 => x"00",
    234 => x"00",
    235 => x"00",
    others => x"00"
    );

begin

    -- Assemble 32-bit instruction from 4 consecutive bytes (little-endian)
    instr_data <= rom_array(to_integer(unsigned(instr_addr) + 3)) &
            rom_array(to_integer(unsigned(instr_addr) + 2)) &
            rom_array(to_integer(unsigned(instr_addr) + 1)) &
            rom_array(to_integer(unsigned(instr_addr)));

    data_data <= rom_array(to_integer(unsigned(data_addr) + 3)) &
            rom_array(to_integer(unsigned(data_addr) + 2)) &
            rom_array(to_integer(unsigned(data_addr) + 1)) &
            rom_array(to_integer(unsigned(data_addr)));

end rom_arch;

