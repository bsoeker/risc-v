library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity rom is
    generic (
        addr_width  : integer := 10  -- 1024 words = 4KB
    );
    port (
        instr_addr : in  std_logic_vector(addr_width + 1 downto 0); -- Byte address (PC)
        instr_data : out std_logic_vector(31 downto 0);  -- Full 32-bit instruction
        data_addr  : in  std_logic_vector(addr_width + 1 downto 0); -- Byte address (ALU)
        data_data  : out std_logic_vector(31 downto 0)  -- Full 32-bit data
    );
end rom;

architecture rom_arch of rom is
    signal instr_word_addr : integer range 0 to 2**addr_width - 1;
    signal data_word_addr  : integer range 0 to 2**addr_width - 1;

    type rom_type is array (0 to 2**addr_width - 1) of std_logic_vector(31 downto 0);
    signal rom_array : rom_type := (
    0 => x"10001117",
    1 => x"00010113",
    2 => x"2E800513",
    3 => x"10000597",
    4 => x"FF458593",
    5 => x"10000617",
    6 => x"FEC60613",
    7 => x"00C58C63",
    8 => x"00054283",
    9 => x"00558023",
    10 => x"00150513",
    11 => x"00158593",
    12 => x"FEDFF06F",
    13 => x"10000517",
    14 => x"FCC50513",
    15 => x"10000597",
    16 => x"FC458593",
    17 => x"00B50863",
    18 => x"00052023",
    19 => x"00450513",
    20 => x"FF5FF06F",
    21 => x"20C000EF",
    22 => x"0000006F",
    23 => x"FE010113",
    24 => x"00112E23",
    25 => x"00812C23",
    26 => x"02010413",
    27 => x"FE042623",
    28 => x"0100006F",
    29 => x"FEC42783",
    30 => x"00178793",
    31 => x"FEF42623",
    32 => x"FEC42703",
    33 => x"000017B7",
    34 => x"9C378793",
    35 => x"FEE7D4E3",
    36 => x"00000013",
    37 => x"00000013",
    38 => x"01C12083",
    39 => x"01812403",
    40 => x"02010113",
    41 => x"00008067",
    42 => x"FE010113",
    43 => x"00112E23",
    44 => x"00812C23",
    45 => x"02010413",
    46 => x"FEA42623",
    47 => x"00000013",
    48 => x"300007B7",
    49 => x"00878793",
    50 => x"0007A783",
    51 => x"0017F793",
    52 => x"FE0788E3",
    53 => x"300007B7",
    54 => x"FEC42703",
    55 => x"00E7A023",
    56 => x"F7DFF0EF",
    57 => x"00000013",
    58 => x"01C12083",
    59 => x"01812403",
    60 => x"02010113",
    61 => x"00008067",
    62 => x"FF010113",
    63 => x"00112623",
    64 => x"00812423",
    65 => x"01010413",
    66 => x"000107B7",
    67 => x"4C078513",
    68 => x"F99FF0EF",
    69 => x"000207B7",
    70 => x"4A878513",
    71 => x"F8DFF0EF",
    72 => x"000307B7",
    73 => x"40078513",
    74 => x"F81FF0EF",
    75 => x"000407B7",
    76 => x"40178513",
    77 => x"F75FF0EF",
    78 => x"00000013",
    79 => x"00C12083",
    80 => x"00812403",
    81 => x"01010113",
    82 => x"00008067",
    83 => x"FF010113",
    84 => x"00112623",
    85 => x"00812423",
    86 => x"01010413",
    87 => x"000507B7",
    88 => x"4FF78513",
    89 => x"F45FF0EF",
    90 => x"000607B7",
    91 => x"4FF78513",
    92 => x"F39FF0EF",
    93 => x"000707B7",
    94 => x"4FF78513",
    95 => x"F2DFF0EF",
    96 => x"000807B7",
    97 => x"40078513",
    98 => x"F21FF0EF",
    99 => x"00000013",
    100 => x"00C12083",
    101 => x"00812403",
    102 => x"01010113",
    103 => x"00008067",
    104 => x"FF010113",
    105 => x"00112623",
    106 => x"00812423",
    107 => x"01010413",
    108 => x"000907B7",
    109 => x"4DE78513",
    110 => x"EF1FF0EF",
    111 => x"000A07B7",
    112 => x"4AD78513",
    113 => x"EE5FF0EF",
    114 => x"000B07B7",
    115 => x"4BE78513",
    116 => x"ED9FF0EF",
    117 => x"000C07B7",
    118 => x"4EF78513",
    119 => x"ECDFF0EF",
    120 => x"000D07B7",
    121 => x"4CA78513",
    122 => x"EC1FF0EF",
    123 => x"000E07B7",
    124 => x"4FE78513",
    125 => x"EB5FF0EF",
    126 => x"00000013",
    127 => x"00C12083",
    128 => x"00812403",
    129 => x"01010113",
    130 => x"00008067",
    131 => x"FF010113",
    132 => x"00112623",
    133 => x"00812423",
    134 => x"01010413",
    135 => x"000F07B7",
    136 => x"4C078513",
    137 => x"E85FF0EF",
    138 => x"001007B7",
    139 => x"4A878513",
    140 => x"E79FF0EF",
    141 => x"001107B7",
    142 => x"40078513",
    143 => x"E6DFF0EF",
    144 => x"001207B7",
    145 => x"40278513",
    146 => x"E61FF0EF",
    147 => x"00000013",
    148 => x"00C12083",
    149 => x"00812403",
    150 => x"01010113",
    151 => x"00008067",
    152 => x"FE010113",
    153 => x"00112E23",
    154 => x"00812C23",
    155 => x"02010413",
    156 => x"FE042623",
    157 => x"0100006F",
    158 => x"FEC42783",
    159 => x"00178793",
    160 => x"FEF42623",
    161 => x"FEC42703",
    162 => x"002627B7",
    163 => x"59F78793",
    164 => x"FEE7D4E3",
    165 => x"E65FF0EF",
    166 => x"EB5FF0EF",
    167 => x"F05FF0EF",
    168 => x"F6DFF0EF",
    169 => x"FE042423",
    170 => x"0100006F",
    171 => x"FE842783",
    172 => x"00178793",
    173 => x"FEF42423",
    174 => x"FE842703",
    175 => x"002627B7",
    176 => x"59F78793",
    177 => x"FEE7D4E3",
    178 => x"00390537",
    179 => x"DDDFF0EF",
    180 => x"00000793",
    181 => x"00078513",
    182 => x"01C12083",
    183 => x"01812403",
    184 => x"02010113",
    185 => x"00008067",
    others => x"00000000"
);

begin
    instr_word_addr <= to_integer(shift_right(unsigned(instr_addr), 2));
    data_word_addr <= to_integer(shift_right(unsigned(data_addr), 2));

    instr_data <= rom_array(instr_word_addr);
    data_data  <= rom_array(data_word_addr);

end rom_arch;

