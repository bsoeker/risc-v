library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity rom is
    generic (
        addr_width  : integer := 10;  -- 2^10 = 1KB
        data_width  : integer := 32 
    );
    port (
        addr : in  std_logic_vector(addr_width - 1 downto 0); -- Byte address (PC)
        data : out std_logic_vector(data_width - 1 downto 0)  -- Full 32-bit instruction
    );
end rom;

architecture rom_arch of rom is

    -- Byte-addressable ROM: Each address holds 1 byte
    type rom_type is array (0 to 2**addr_width - 1) of std_logic_vector(7 downto 0);
    signal rom_array : rom_type := (
    0 => x"17",
    1 => x"11",
    2 => x"00",
    3 => x"10",
    4 => x"13",
    5 => x"01",
    6 => x"01",
    7 => x"00",
    8 => x"13",
    9 => x"05",
    10 => x"40",
    11 => x"0B",
    12 => x"97",
    13 => x"05",
    14 => x"00",
    15 => x"10",
    16 => x"93",
    17 => x"85",
    18 => x"45",
    19 => x"FF",
    20 => x"17",
    21 => x"06",
    22 => x"00",
    23 => x"10",
    24 => x"13",
    25 => x"06",
    26 => x"26",
    27 => x"FF",
    28 => x"63",
    29 => x"8C",
    30 => x"C5",
    31 => x"00",
    32 => x"83",
    33 => x"42",
    34 => x"05",
    35 => x"00",
    36 => x"23",
    37 => x"80",
    38 => x"55",
    39 => x"00",
    40 => x"13",
    41 => x"05",
    42 => x"15",
    43 => x"00",
    44 => x"93",
    45 => x"85",
    46 => x"15",
    47 => x"00",
    48 => x"6F",
    49 => x"F0",
    50 => x"DF",
    51 => x"FE",
    52 => x"17",
    53 => x"05",
    54 => x"00",
    55 => x"10",
    56 => x"13",
    57 => x"05",
    58 => x"25",
    59 => x"FD",
    60 => x"97",
    61 => x"05",
    62 => x"00",
    63 => x"10",
    64 => x"93",
    65 => x"85",
    66 => x"A5",
    67 => x"FC",
    68 => x"63",
    69 => x"08",
    70 => x"B5",
    71 => x"00",
    72 => x"23",
    73 => x"20",
    74 => x"05",
    75 => x"00",
    76 => x"13",
    77 => x"05",
    78 => x"45",
    79 => x"00",
    80 => x"6F",
    81 => x"F0",
    82 => x"5F",
    83 => x"FF",
    84 => x"EF",
    85 => x"00",
    86 => x"80",
    87 => x"00",
    88 => x"6F",
    89 => x"00",
    90 => x"00",
    91 => x"00",
    92 => x"13",
    93 => x"01",
    94 => x"01",
    95 => x"FE",
    96 => x"23",
    97 => x"2E",
    98 => x"11",
    99 => x"00",
    100 => x"23",
    101 => x"2C",
    102 => x"81",
    103 => x"00",
    104 => x"13",
    105 => x"04",
    106 => x"01",
    107 => x"02",
    108 => x"B7",
    109 => x"07",
    110 => x"00",
    111 => x"20",
    112 => x"93",
    113 => x"87",
    114 => x"47",
    115 => x"00",
    116 => x"83",
    117 => x"A7",
    118 => x"07",
    119 => x"00",
    120 => x"93",
    121 => x"F7",
    122 => x"17",
    123 => x"00",
    124 => x"23",
    125 => x"26",
    126 => x"F4",
    127 => x"FE",
    128 => x"83",
    129 => x"27",
    130 => x"C4",
    131 => x"FE",
    132 => x"93",
    133 => x"F7",
    134 => x"F7",
    135 => x"0F",
    136 => x"93",
    137 => x"87",
    138 => x"17",
    139 => x"04",
    140 => x"A3",
    141 => x"05",
    142 => x"F4",
    143 => x"FE",
    144 => x"B7",
    145 => x"07",
    146 => x"00",
    147 => x"20",
    148 => x"03",
    149 => x"47",
    150 => x"B4",
    151 => x"FE",
    152 => x"23",
    153 => x"A0",
    154 => x"E7",
    155 => x"00",
    156 => x"93",
    157 => x"07",
    158 => x"00",
    159 => x"00",
    160 => x"13",
    161 => x"85",
    162 => x"07",
    163 => x"00",
    164 => x"83",
    165 => x"20",
    166 => x"C1",
    167 => x"01",
    168 => x"03",
    169 => x"24",
    170 => x"81",
    171 => x"01",
    172 => x"13",
    173 => x"01",
    174 => x"01",
    175 => x"02",
    176 => x"67",
    177 => x"80",
    178 => x"00",
    179 => x"00",
    180 => x"48",
    181 => x"65",
    182 => x"6C",
    183 => x"6C",
    184 => x"6F",
    185 => x"00",
    186 => x"00",
    187 => x"00",
    others => x"00"
    );

begin

    -- Assemble 32-bit instruction from 4 consecutive bytes (little-endian)
    data <= rom_array(to_integer(unsigned(addr) + 3)) &
            rom_array(to_integer(unsigned(addr) + 2)) &
            rom_array(to_integer(unsigned(addr) + 1)) &
            rom_array(to_integer(unsigned(addr)));

end rom_arch;

